// scr1_pkg.sv
package scr1_pkg;
//	`include "scr1_arch_description.svh"
	`include "scr1_riscv_isa_decoding.svh"
endpackage
